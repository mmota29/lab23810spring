library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_mux32to1_32bit is
end tb_mux32to1_32bit;

architecture sim of tb_mux32to1_32bit is
  component mux32to1_32bit
    port(
      i_D : in std_logic_vector(1023 downto 0);
      i_S : in std_logic_vector(4 downto 0);
      o_Y : out std_logic_vector(31 downto 0)
    );
  end component;

  signal d : std_logic_vector(1023 downto 0) := (others => '0');
  signal s : std_logic_vector(4 downto 0) := (others => '0');
  signal y : std_logic_vector(31 downto 0);

  procedure set_word(signal big : inout std_logic_vector(1023 downto 0); idx : integer; val : std_logic_vector(31 downto 0)) is
  begin
    big((idx*32 + 31) downto (idx*32)) <= val;
  end procedure;

begin
  uut: mux32to1_32bit
    port map(
      i_D => d,
      i_S => s,
      o_Y => y
    );

  stim: process
  begin
    -- fill with 0..31
    for i in 0 to 31 loop
      set_word(d, i, std_logic_vector(to_unsigned(i, 32)));
    end loop;

    s <= "00000"; wait for 10 ns; -- expect 0
    s <= "00001"; wait for 10 ns; -- expect 1
    s <= "01001"; wait for 10 ns; -- expect 9
    s <= "11111"; wait for 10 ns; -- expect 31

    -- change these
    set_word(d, 5, x"4D494348"); -- "MICH"
    set_word(d, 6, x"41454C00"); -- "AEL\0"
    s <= "00101"; wait for 10 ns;
    s <= "00110"; wait for 10 ns;

    wait;
  end process;
end sim;