    Mac OS X            	   2  >     p    ��������                          ATTR      p   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     4   <  com.apple.quarantine M��h    �׳     @6�02�I����T;�J                                                      q/0281;69710905;Chrome;EA1CF270-A450-475B-8D21-B9BA413E4C34 