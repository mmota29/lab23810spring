    Mac OS X            	   2   �      �    ��������                          ATTR       �   �   <                  �   <  com.apple.quarantine q/0281;69710905;Chrome;EA1CF270-A450-475B-8D21-B9BA413E4C34 